<!doctype html public "-//W3C//DTD HTML 3.2 Final//EN">
<html>
 <head>
  <title>Testsida f&ouml;r Apache-installationen</title>
 </head>
<!-- Background white, links blue (unvisited), navy (visited), red (active) -->
 <body
  bgcolor="#FFFFFF"
  text="#000000"
  link="#0000FF"
  vlink="#000080"
  alink="#FF0000"
 >
  <h1 align="CENTER">
   Det fungerade! Apache &auml;r installerad p&aring; denna maskin!
  </h1>
  <p>
  Om du kan se denna sida s&aring; har &auml;garen till denna maskin installerat
  webbserverprogramvaran Apache.<br>
  Denne m&aring;ste nu placera webbsidor i detta bibliotek och &auml;ndra p&aring; denna sida, eller
  peka servern mot ett annat bibliotek.
  </p>
  <hr>
  <blockquote>
   Om du f&ouml;rv&auml;ntat dig att se n&aring;got helt annat h&auml;r &auml;n denna sida, <strong>kontakta
   v&auml;nligen administrat&ouml;ren f&ouml;r den webbserver du f&ouml;rs&ouml;ker komma i kontakt med.</strong>
   (F&ouml;rs&ouml;k att skicka ett brev till <samp>&lt;webmaster@<em>domain</em>&gt;</samp>.)
   Apache Software Foundation har inget med denna webbplats att g&ouml;ra, s&aring; det &auml;r ingen id&eacute;
   att skicka mail till f&ouml;rfattarna av Apache r&ouml;rande denna webbplats.
  </blockquote>
  <hr>
  <p>
  Apache-<a href="manual/">dokumentationen</a> &auml;r inkluderad i denna distribution.
  </p>
  <p>
  Administrat&ouml;ren av denna webbplats f&aring;r g&auml;rna anv&auml;nda f&ouml;ljande bild till en webbplats som anv&auml;nder Apache.<br>
  Tack f&ouml;r att ni anv&auml;nder Apache!
  </p>
  <div align="CENTER">
   <img src="apache_pb.gif" alt="">
  </div>
 </body>
</html>
